module Top (
	input i_rst_n,
	input i_clk,
	input i_key_0,			
	input i_key_1,			
	input i_key_2,			
	input [2:0] i_speed,	
	input i_fast,			
	input i_slow_0, 
	input i_slow_1,
	input	i_reverse,	
	
	// AudDSP and SRAM
	output [19:0] o_SRAM_ADDR,
	inout  [15:0] io_SRAM_DQ,
	output        o_SRAM_WE_N,
	output        o_SRAM_CE_N,
	output        o_SRAM_OE_N,
	output        o_SRAM_LB_N,
	output        o_SRAM_UB_N,
	
	// I2C
	input  i_clk_100k,
	output o_I2C_SCLK,
	inout  io_I2C_SDAT,
	
	// AudPlayer
	input  i_AUD_ADCDAT,
	inout  i_AUD_ADCLRCK,
	inout  i_AUD_BCLK,
	inout  i_AUD_DACLRCK,
	output o_AUD_DACDAT,
	
	output [3:0] o_state,
	//output [2:0] o_voice_state,

	// SEVENDECODER (optional display)
	// output [5:0] o_record_time,
	// output [5:0] o_play_time,

	// LCD (optional display)
	// input        i_clk_800k,
	// inout  [7:0] o_LCD_DATA,
	// output       o_LCD_EN,
	// output       o_LCD_RS,
	// output       o_LCD_RW,
	// output       o_LCD_ON,
	// output       o_LCD_BLON,

	// LED
	// output  [8:0] o_ledg,
	//output [17:0] o_led,
	output o_vol,
	output o_volume
);

// design the FSM and states as you like
parameter S_IDLE       = 0;
parameter S_I2CED      = 1;
parameter S_RECD       = 2;
parameter S_RECD_PAUSE = 3;
parameter S_PLAY       = 4;
parameter S_PLAY_PAUSE = 5;

logic [3:0] state_w, state_r;
logic i2c_oen, i2c_sdat;
logic [19:0] addr_record, addr_play, end_addr_r, end_addr_w;
logic [15:0] data_record, data_play, dac_data;

//logic [3:0] recent_state_w, recent_state_r;


assign io_I2C_SDAT = (i2c_oen) ? i2c_sdat : 1'bz;

assign o_SRAM_ADDR = (state_r == S_RECD || state_r == S_RECD_PAUSE) ? addr_record : addr_play[19:0];
assign io_SRAM_DQ  = (state_r == S_RECD || state_r == S_RECD_PAUSE) ? data_record : 16'dz; // sram_dq as output
assign data_play   = (state_r == S_RECD || state_r == S_RECD_PAUSE) ? 16'd0 : io_SRAM_DQ; // sram_dq as input

assign o_SRAM_WE_N = (state_r==S_RECD || state_r == S_RECD_PAUSE) ? 1'b0 : 1'b1;
assign o_SRAM_CE_N = 1'b0;
assign o_SRAM_OE_N = 1'b0;
assign o_SRAM_LB_N = 1'b0;
assign o_SRAM_UB_N = 1'b0;
logic i2c_finish;
assign o_state = state_r;



// below is a simple example for module division
// you can design these as you like

// === I2cInitializer ===
// sequentially sent out settings to initialize WM8731 with I2C protocal

I2CInitializer init0(
	.i_rst_n(i_rst_n),
	.i_clk(i_clk_100k),
	.i_start(1),
	.o_finished(i2c_finish),
	.o_sclk(o_I2C_SCLK),
	.o_sdat(i2c_sdat),
	.o_oen(i2c_oen) // you are outputing (you are not outputing only when you are "ack"ing.)
);

// === AudDSP ===
// responsible for DSP operations including fast play and slow play at different speed
// in other words, determine which data addr to be fetch for player 
logic audplayer_en;
AudDSP dsp0(
	.i_rst_n(i_rst_n),
	.i_clk(i_clk),
	.i_start(state_r==S_PLAY),
	.i_pause(state_r==S_PLAY_PAUSE),
	.i_stop(state_r==S_I2CED),
	.i_speed(i_speed),
	.i_fast(i_fast),
	.i_slow_0(i_slow_0), // constant interpolation
	.i_slow_1(i_slow_1), // linear interpolation
	.i_reverse(i_reverse),
	.i_daclrck(i_AUD_DACLRCK),
	.i_sram_data(data_play),
	.i_end_address(end_addr_w),
	.o_dac_data(dac_data),
	.o_sram_addr(addr_play),
	.o_audplayer_en(audplayer_en)
);

// === AudPlayer ===
// receive data address from DSP and fetch data to sent to WM8731 with I2S protocal
AudPlayer player0(
	.i_rst_n(i_rst_n),
	.i_bclk(i_AUD_BCLK),
	.i_daclrck(i_AUD_DACLRCK),
	.i_en(audplayer_en), // enable AudPlayer only when playing audio, work with AudDSP
	.i_dac_data(dac_data), //dac_data
	.o_aud_dacdat(o_AUD_DACDAT)
);

// === AudRecorder ===
// receive data from WM8731 with I2S protocal and save to SRAM
AudRecorder recorder0(
	.i_rst_n(i_rst_n), 
	.i_clk(i_AUD_BCLK),
	.i_lrc(i_AUD_ADCLRCK),
	.i_start(state_r==S_RECD),
	.i_pause(state_r==S_RECD_PAUSE),
	.i_stop(state_r==S_I2CED),
	.i_data(i_AUD_ADCDAT),
	.o_address(addr_record),
	.o_data(data_record)
);
Volume volume(
	.i_rst_n(i_rst_n), 
	.i_clk(i_AUD_BCLK),
	.i_data(data_record),
	.i_recording(state_r==S_RECD),
	//.o_state(o_voice_state),
	//.o_led(o_led),
	.o_vol(o_vol),
	.o_volume(o_volume)
);

always_comb begin
	// design your control here
	state_w = state_r;
	//recent_state_w = recent_state_r;
	end_addr_w = end_addr_r;
	case(state_r) 
		S_IDLE: begin
			state_w = (i2c_finish)? S_I2CED : state_r;
		end
		S_I2CED: begin
			
			if(i_key_0) begin
				state_w = S_RECD;
			end 
			else if(i_key_1) begin
				state_w = S_PLAY;
			end
		end
		S_RECD: begin
			if(i_key_0) begin
				state_w = S_RECD_PAUSE;
			end
			else if(i_key_2) begin
				state_w = S_I2CED;
				end_addr_w = addr_record;
			end
			
		end
		
		S_RECD_PAUSE: begin
			if(i_key_0) begin
				state_w = S_RECD;
			end
			else if(i_key_2) begin
				state_w = S_I2CED;
				end_addr_w = addr_record;
			end

		end
		S_PLAY: begin
			if(i_key_1) begin
				state_w = S_PLAY_PAUSE;
			end
			else if(i_key_2) begin
				state_w = S_I2CED;
			end
			
		end
		S_PLAY_PAUSE: begin
			if(i_key_1) begin
				state_w = S_PLAY;
			end
			else if(i_key_2) begin
				state_w = S_I2CED;
			end

		end
	endcase	



end

always_ff @(posedge i_AUD_BCLK or negedge i_rst_n) begin
	if (!i_rst_n) begin
		state_r <= S_IDLE;
		end_addr_r <= 20'b0;
		
	end
	else begin
		state_r <= state_w;
		end_addr_r <= end_addr_w;
		
	end
end

endmodule